library ieee;
use ieee.std_logic_1164.all;

library work;
use work.font.all;

package font_4x6 is

  constant font_4x6_c : font_t :=
    font_define(
      4, 6,
      glyph( -- '^@' 0x00
        "    ",
        "    ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '^A' 0x01
        " ## ",
        "#  #",
        "#  #",
        "####",
        " ## ",
        "    ") &
      glyph( -- '^B' 0x02
        " ## ",
        "####",
        "####",
        "#  #",
        " ## ",
        "    ") &
      glyph( -- '^C' 0x03
        "    ",
        "# # ",
        "### ",
        "### ",
        " #  ",
        "    ") &
      glyph( -- '^D' 0x04
        "    ",
        " #  ",
        "### ",
        " #  ",
        "    ",
        "    ") &
      glyph( -- '^E' 0x05
        "    ",
        " #  ",
        "# # ",
        " #  ",
        "### ",
        "    ") &
      glyph( -- '^F' 0x06
        "    ",
        " #  ",
        "### ",
        " #  ",
        "### ",
        "    ") &
      glyph( -- '^G' 0x07
        "    ",
        "    ",
        " ## ",
        " ## ",
        "    ",
        "    ") &
      glyph( -- '^H' 0x08
        "####",
        "####",
        "#  #",
        "#  #",
        "####",
        "####") &
      glyph( -- '^I' 0x09
        "    ",
        " ## ",
        "#  #",
        " ## ",
        "    ",
        "    ") &
      glyph( -- '^J' 0x0A
        "####",
        "#  #",
        " ## ",
        "#  #",
        "####",
        "####") &
      glyph( -- '^K' 0x0B
        " ###",
        "  ##",
        " #  ",
        "# ##",
        " ## ",
        "    ") &
      glyph( -- '^L' 0x0C
        " ## ",
        "#  #",
        " ## ",
        "  # ",
        " ###",
        "  # ") &
      glyph( -- '^M' 0x0D
        "  # ",
        "  ##",
        "  # ",
        "  # ",
        "##  ",
        "##  ") &
      glyph( -- '^N' 0x0E
        " ###",
        " # #",
        " # #",
        " # #",
        "## #",
        "## #") &
      glyph( -- '^O' 0x0F
        "# # ",
        " ###",
        " # #",
        " ## ",
        " # #",
        "    ") &
      glyph( -- '^P' 0x10
        "#   ",
        "##  ",
        "### ",
        "##  ",
        "#   ",
        "    ") &
      glyph( -- '^Q' 0x11
        "  # ",
        " ## ",
        "### ",
        " ## ",
        "  # ",
        "    ") &
      glyph( -- '^R' 0x12
        " #  ",
        "### ",
        " #  ",
        "### ",
        " #  ",
        "    ") &
      glyph( -- '^S' 0x13
        "# # ",
        "# # ",
        "# # ",
        "    ",
        "# # ",
        "    ") &
      glyph( -- '^T' 0x14
        " ###",
        "# ##",
        " ###",
        "  ##",
        "  ##",
        "    ") &
      glyph( -- '^U' 0x15
        " ###",
        "##  ",
        "### ",
        " ## ",
        "##  ",
        "    ") &
      glyph( -- '^V' 0x16
        "    ",
        "    ",
        "    ",
        "### ",
        "### ",
        "    ") &
      glyph( -- '^W' 0x17
        " #  ",
        "### ",
        " #  ",
        "### ",
        " #  ",
        "####") &
      glyph( -- '^X' 0x18
        " #  ",
        "### ",
        " #  ",
        " #  ",
        " #  ",
        "    ") &
      glyph( -- '^Y' 0x19
        " #  ",
        " #  ",
        " #  ",
        "### ",
        " #  ",
        "    ") &
      glyph( -- '^Z' 0x1A
        " #  ",
        "  # ",
        "####",
        "  # ",
        " #  ",
        "    ") &
      glyph( -- '^[' 0x1B
        "  # ",
        " #  ",
        "####",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '^\' 0x1C
        "    ",
        "    ",
        "#   ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- '^]' 0x1D
        "    ",
        "#  #",
        "####",
        "#  #",
        "    ",
        "    ") &
      glyph( -- '^^' 0x1E
        "    ",
        " #  ",
        " ## ",
        "### ",
        "####",
        "    ") &
      glyph( -- '^_' 0x1F
        "    ",
        "####",
        "### ",
        " ## ",
        " #  ",
        "    ") &
      glyph( -- ' ' 0x20
        "    ",
        "    ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '!' 0x21
        " #  ",
        " #  ",
        " #  ",
        "    ",
        " #  ",
        "    ") &
      glyph( -- '"' 0x22
        "# # ",
        "# # ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '#' 0x23
        "# # ",
        "### ",
        "# # ",
        "### ",
        "# # ",
        "    ") &
      glyph( -- '$' 0x24
        " ## ",
        "##  ",
        "### ",
        " ## ",
        "##  ",
        "    ") &
      glyph( -- '%' 0x25
        "# # ",
        "  # ",
        " #  ",
        "#   ",
        "# # ",
        "    ") &
      glyph( -- '&' 0x26
        " ## ",
        "# # ",
        " # #",
        "# # ",
        "## #",
        "    ") &
      glyph( -- ''' 0x27
        " #  ",
        " #  ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '(' 0x28
        " #  ",
        "#   ",
        "#   ",
        "#   ",
        " #  ",
        "    ") &
      glyph( -- ')' 0x29
        " #  ",
        "  # ",
        "  # ",
        "  # ",
        " #  ",
        "    ") &
      glyph( -- '*' 0x2A
        "# # ",
        " #  ",
        "### ",
        " #  ",
        "# # ",
        "    ") &
      glyph( -- '+' 0x2B
        "    ",
        " #  ",
        "### ",
        " #  ",
        "    ",
        "    ") &
      glyph( -- ',' 0x2C
        "    ",
        "    ",
        "    ",
        "    ",
        " #  ",
        "#   ") &
      glyph( -- '-' 0x2D
        "    ",
        "    ",
        "### ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '.' 0x2E
        "    ",
        "    ",
        "    ",
        "    ",
        " #  ",
        "    ") &
      glyph( -- '/' 0x2F
        "  # ",
        " #  ",
        " #  ",
        " #  ",
        "#   ",
        "    ") &
      glyph( -- '0' 0x30
        " ## ",
        "# # ",
        "# # ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- '1' 0x31
        " #  ",
        "##  ",
        " #  ",
        " #  ",
        "### ",
        "    ") &
      glyph( -- '2' 0x32
        " ## ",
        "# # ",
        "  # ",
        " # ",
        "### ",
        "    ") &
      glyph( -- '3' 0x33
        "### ",
        "  # ",
        " #  ",
        "  # ",
        "##  ",
        "    ") &
      glyph( -- '4' 0x34
        "  # ",
        " ## ",
        "# # ",
        "####",
        "  # ",
        "    ") &
      glyph( -- '5' 0x35
        "### ",
        "#   ",
        "##  ",
        "  # ",
        "##  ",
        "    ") &
      glyph( -- '6' 0x36
        " ## ",
        "#   ",
        "### ",
        "#  #",
        " ## ",
        "    ") &
      glyph( -- '7' 0x37
        "### ",
        "  # ",
        " #  ",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- '8' 0x38
        " ## ",
        "# # ",
        " #  ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- '9' 0x39
        " ## ",
        "# # ",
        " ## ",
        "  # ",
        "##  ",
        "    ") &
      glyph( -- ':' 0x3A
        "    ",
        " #  ",
        "    ",
        " #  ",
        "    ",
        "    ") &
      glyph( -- ';' 0x3B
        "    ",
        "    ",
        " #  ",
        "    ",
        " #  ",
        "#   ") &
      glyph( -- '<' 0x3C
        "  # ",
        " #  ",
        "#   ",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '=' 0x3D
        "    ",
        "### ",
        "    ",
        "### ",
        "    ",
        "    ") &
      glyph( -- '>' 0x3E
        "#   ",
        " #  ",
        "  # ",
        " #  ",
        "#   ",
        "    ") &
      glyph( -- '?' 0x3F
        "##  ",
        "  # ",
        " #  ",
        "    ",
        " #  ",
        "    ") &
      glyph( -- '@' 0x40
        " #  ",
        "# # ",
        "# # ",
        "#   ",
        " ## ",
        "    ") &
      glyph( -- 'A' 0x41
        " ## ",
        "# # ",
        "### ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'B' 0x42
        "##  ",
        "# # ",
        "##  ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'C' 0x43
        " ## ",
        "#   ",
        "#   ",
        "#   ",
        " ## ",
        "    ") &
      glyph( -- 'D' 0x44
        "##  ",
        "# # ",
        "# # ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'E' 0x45
        " ## ",
        "#   ",
        "##  ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- 'F' 0x46
        " ## ",
        "#   ",
        "### ",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- 'G' 0x47
        " ## ",
        "#   ",
        "# # ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'H' 0x48
        "# # ",
        "# # ",
        "### ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'I' 0x49
        "### ",
        " #  ",
        " #  ",
        " #  ",
        "### ",
        "    ") &
      glyph( -- 'J' 0x4A
        "### ",
        "  # ",
        "  # ",
        "  # ",
        "##  ",
        "    ") &
      glyph( -- 'K' 0x4B
        "#   ",
        "# # ",
        "##  ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'L' 0x4C
        "#   ",
        "#   ",
        "#   ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- 'M' 0x4D
        " ## ",
        "### ",
        "# # ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'N' 0x4E
        "##  ",
        "# # ",
        "# # ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'O' 0x4F
        " ## ",
        "# # ",
        "# # ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'P' 0x50
        "##  ",
        "# # ",
        "##  ",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- 'Q' 0x51
        " ## ",
        "# # ",
        "# # ",
        "# # ",
        "### ",
        "    ") &
      glyph( -- 'R' 0x52
        "##  ",
        "# # ",
        "##  ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'S' 0x53
        " ## ",
        "#   ",
        " #  ",
        "  # ",
        "##  ",
        "    ") &
      glyph( -- 'T' 0x54
        "### ",
        " #  ",
        " #  ",
        " #  ",
        " #  ",
        "    ") &
      glyph( -- 'U' 0x55
        "# # ",
        "# # ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- 'V' 0x56
        "# # ",
        "# # ",
        "# # ",
        "# # ",
        " #  ",
        "    ") &
      glyph( -- 'W' 0x57
        "# # ",
        "# # ",
        "### ",
        "### ",
        "# # ",
        "    ") &
      glyph( -- 'X' 0x58
        "# # ",
        "# # ",
        " #  ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'Y' 0x59
        "# # ",
        "# # ",
        " #  ",
        " #  ",
        " #  ",
        "    ") &
      glyph( -- 'Z' 0x5A
        "### ",
        "  # ",
        " #  ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- '[' 0x5B
        "##  ",
        "#   ",
        "#   ",
        "#   ",
        "##  ",
        "    ") &
      glyph( -- '\' 0x5C
        "#   ",
        "#   ",
        " #  ",
        "  # ",
        "  # ",
        "    ") &
      glyph( -- ']' 0x5D
        " ## ",
        "  # ",
        "  # ",
        "  # ",
        " ## ",
        "    ") &
      glyph( -- '^' 0x5E
        " #  ",
        "# # ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '_' 0x5F
        "    ",
        "    ",
        "    ",
        "    ",
        "    ",
        "####") &
      glyph( -- '`' 0x60
        "#   ",
        " #  ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- 'a' 0x61
        "    ",
        "    ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- 'b' 0x62
        "#   ",
        "#   ",
        "##  ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'c' 0x63
        "    ",
        "    ",
        " ## ",
        "#   ",
        " ## ",
        "    ") &
      glyph( -- 'd' 0x64
        "  # ",
        "  # ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- 'e' 0x65
        "    ",
        "    ",
        "### ",
        "##  ",
        " ## ",
        "    ") &
      glyph( -- 'f' 0x66
        " ## ",
        "#   ",
        "##  ",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- 'g' 0x67
        "    ",
        "    ",
        " ## ",
        "### ",
        "  # ",
        "##  ") &
      glyph( -- 'h' 0x68
        "#   ",
        "#   ",
        "##  ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'i' 0x69
        " #  ",
        "    ",
        " #  ",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- 'j' 0x6A
        " #  ",
        "    ",
        " #  ",
        " #  ",
        " #  ",
        "#   ") &
      glyph( -- 'k' 0x6B
        "#   ",
        "#   ",
        "# # ",
        "##  ",
        "# # ",
        "    ") &
      glyph( -- 'l' 0x6C
        "#   ",
        "#   ",
        "#   ",
        "#   ",
        " #  ",
        "    ") &
      glyph( -- 'm' 0x6D
        "    ",
        "    ",
        "##  ",
        "### ",
        "# # ",
        "    ") &
      glyph( -- 'n' 0x6E
        "    ",
        "    ",
        "##  ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- 'o' 0x6F
        "    ",
        "    ",
        " ## ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'p' 0x70
        "    ",
        "    ",
        "##  ",
        "# # ",
        "##  ",
        "#   ") &
      glyph( -- 'q' 0x71
        "    ",
        "    ",
        " ## ",
        "# # ",
        " ## ",
        "  # ") &
      glyph( -- 'r' 0x72
        "    ",
        "    ",
        " ## ",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- 's' 0x73
        "    ",
        "    ",
        " ## ",
        " #  ",
        "##  ",
        "    ") &
      glyph( -- 't' 0x74
        "#   ",
        "##  ",
        "#   ",
        "#   ",
        " #  ",
        "    ") &
      glyph( -- 'u' 0x75
        "    ",
        "    ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- 'v' 0x76
        "    ",
        "    ",
        "# # ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- 'w' 0x77
        "    ",
        "    ",
        "# # ",
        "### ",
        "##  ",
        "    ") &
      glyph( -- 'x' 0x78
        "    ",
        "    ",
        "# # ",
        " #  ",
        "# # ",
        "    ") &
      glyph( -- 'y' 0x79
        "    ",
        "    ",
        "# # ",
        " ## ",
        "  # ",
        "##  ") &
      glyph( -- 'z' 0x7A
        "    ",
        "    ",
        "### ",
        " #  ",
        "  # ",
        "##  ") &
      glyph( -- '{' 0x7B
        " ## ",
        " #  ",
        "#   ",
        " #  ",
        " ## ",
        "    ") &
      glyph( -- '|' 0x7C
        " #  ",
        " #  ",
        " #  ",
        " #  ",
        " #  ",
        "    ") &
      glyph( -- '}' 0x7D
        "##  ",
        " #  ",
        "  # ",
        " #  ",
        "##  ",
        "    ") &
      glyph( -- '~' 0x7E
        "    ",
        " # #",
        "# # ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '' 0x7F
        "    ",
        " #  ",
        "# # ",
        "# # ",
        "### ",
        "    ") &
      glyph( -- '\200' 0x80
        "    ",
        " ## ",
        "#   ",
        " ## ",
        " #  ",
        "#   ") &
      glyph( -- '\201' 0x81
        "# # ",
        "    ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\202' 0x82
        "# # ",
        "    ",
        "### ",
        "##  ",
        " ## ",
        "    ") &
      glyph( -- '\203' 0x83
        " ## ",
        "    ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\204' 0x84
        "# # ",
        "    ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\205' 0x85
        "##  ",
        "    ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\206' 0x86
        "### ",
        " #  ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\207' 0x87
        "    ",
        "    ",
        " ## ",
        "#   ",
        " ## ",
        " #  ") &
      glyph( -- '\210' 0x88
        " ## ",
        "    ",
        "### ",
        "##  ",
        " ## ",
        "    ") &
      glyph( -- '\211' 0x89
        "# # ",
        "    ",
        "### ",
        "##  ",
        " ## ",
        "    ") &
      glyph( -- '\212' 0x8A
        "##  ",
        "    ",
        "### ",
        "##  ",
        " ## ",
        "    ") &
      glyph( -- '\213' 0x8B
        "# # ",
        "    ",
        " #  ",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '\214' 0x8C
        " ## ",
        "    ",
        " #  ",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '\215' 0x8D
        " ## ",
        "    ",
        " #  ",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '\216' 0x8E
        "# # ",
        " #  ",
        "# # ",
        "### ",
        "# # ",
        "    ") &
      glyph( -- '\217' 0x8F
        " #  ",
        " #  ",
        "# # ",
        "### ",
        "# # ",
        "    ") &
      glyph( -- '\220' 0x90
        " #  ",
        "### ",
        "##  ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- '\221' 0x91
        "    ",
        "    ",
        " ## ",
        "# ##",
        " ###",
        "    ") &
      glyph( -- '\222' 0x92
        " ###",
        "# # ",
        "####",
        "# # ",
        "# ##",
        "    ") &
      glyph( -- '\223' 0x93
        " ## ",
        "    ",
        "##  ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\224' 0x94
        "# # ",
        "    ",
        "##  ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\225' 0x95
        " ## ",
        "    ",
        "##  ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\226' 0x96
        " #  ",
        "    ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\227' 0x97
        "#   ",
        " #  ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\230' 0x98
        "# # ",
        "    ",
        "# # ",
        " ## ",
        "  # ",
        "##  ") &
      glyph( -- '\231' 0x99
        "# # ",
        "##  ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\232' 0x9A
        "# # ",
        "    ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\233' 0x9B
        "    ",
        " #  ",
        " ## ",
        "##  ",
        " ## ",
        " #  ") &
      glyph( -- '\234' 0x9C
        " ## ",
        "#   ",
        "##  ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- '\235' 0x9D
        "# # ",
        "# # ",
        " #  ",
        "### ",
        " #  ",
        "    ") &
      glyph( -- '\236' 0x9E
        "##  ",
        "# # ",
        "##  ",
        "# ##",
        "# ##",
        "    ") &
      glyph( -- '\237' 0x9F
        "  # ",
        " #  ",
        "### ",
        " #  ",
        "#   ",
        "    ") &
      glyph( -- '\240' 0xA0
        " ## ",
        "    ",
        " ## ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\241' 0xA1
        " ## ",
        "    ",
        " #  ",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '\242' 0xA2
        " ## ",
        "    ",
        "##  ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\243' 0xA3
        "  # ",
        "    ",
        "# # ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\244' 0xA4
        " # #",
        "  # ",
        "##  ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- '\245' 0xA5
        "  # ",
        "##  ",
        "# # ",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- '\246' 0xA6
        " ## ",
        "# # ",
        " ## ",
        "    ",
        "### ",
        "    ") &
      glyph( -- '\247' 0xA7
        "##  ",
        "# # ",
        " ## ",
        "    ",
        "### ",
        "    ") &
      glyph( -- '\250' 0xA8
        " #  ",
        "    ",
        " #  ",
        "#   ",
        " ## ",
        "    ") &
      glyph( -- '\251' 0xA9
        "    ",
        "    ",
        "####",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- '\252' 0xAA
        "    ",
        "    ",
        "####",
        "   #",
        "   #",
        "    ") &
      glyph( -- '\253' 0xAB
        "#  #",
        "  # ",
        " ## ",
        "#  #",
        "  # ",
        "  ##") &
      glyph( -- '\254' 0xAC
        "#  #",
        "  # ",
        " #  ",
        "# # ",
        " ###",
        "   #") &
      glyph( -- '\255' 0xAD
        " #  ",
        "    ",
        " #  ",
        " #  ",
        " #  ",
        "    ") &
      glyph( -- '\256' 0xAE
        "    ",
        " # #",
        "# # ",
        "# # ",
        " # #",
        "    ") &
      glyph( -- '\257' 0xAF
        "    ",
        "# # ",
        " # #",
        " # #",
        "# # ",
        "    ") &
      glyph( -- '\260' 0xB0
        "  # ",
        "#   ",
        "  # ",
        "#   ",
        "  # ",
        "#   ") &
      glyph( -- '\261' 0xB1
        " # #",
        "# # ",
        " # #",
        "# # ",
        " # #",
        "# # ") &
      glyph( -- '\262' 0xB2
        " ###",
        "## #",
        " ###",
        "## #",
        " ###",
        "## #") &
      glyph( -- '\263' 0xB3
        "  # ",
        "  # ",
        "  # ",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\264' 0xB4
        "  # ",
        "  # ",
        "### ",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\265' 0xB5
        "  # ",
        "  # ",
        "### ",
        "### ",
        "  # ",
        "  # ") &
      glyph( -- '\266' 0xB6
        " ## ",
        " ## ",
        "### ",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\267' 0xB7
        "    ",
        "    ",
        "### ",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\270' 0xB8
        "    ",
        "    ",
        "### ",
        "### ",
        "  # ",
        "  # ") &
      glyph( -- '\271' 0xB9
        " ## ",
        " ## ",
        "### ",
        "### ",
        " ## ",
        " ## ") &
      glyph( -- '\272' 0xBA
        " ## ",
        " ## ",
        " ## ",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\273' 0xBB
        "    ",
        "    ",
        "### ",
        "### ",
        " ## ",
        " ## ") &
      glyph( -- '\274' 0xBC
        " ## ",
        " ## ",
        "### ",
        "### ",
        "    ",
        "    ") &
      glyph( -- '\275' 0xBD
        " ## ",
        " ## ",
        "### ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\276' 0xBE
        "  # ",
        "  # ",
        "### ",
        "### ",
        "    ",
        "    ") &
      glyph( -- '\277' 0xBF
        "    ",
        "    ",
        "### ",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\300' 0xC0
        "  # ",
        "  # ",
        "  ##",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\301' 0xC1
        "  # ",
        "  # ",
        "####",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\302' 0xC2
        "    ",
        "    ",
        "####",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\303' 0xC3
        "  # ",
        "  # ",
        "  ##",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\304' 0xC4
        "    ",
        "    ",
        "####",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\305' 0xC5
        "  # ",
        "  # ",
        "####",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\306' 0xC6
        "  # ",
        "  # ",
        "  ##",
        "  ##",
        "  # ",
        "  # ") &
      glyph( -- '\307' 0xC7
        " ## ",
        " ## ",
        " ###",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\310' 0xC8
        " ## ",
        " ## ",
        " ###",
        " ###",
        "    ",
        "    ") &
      glyph( -- '\311' 0xC9
        "    ",
        "    ",
        " ###",
        " ###",
        " ## ",
        " ## ") &
      glyph( -- '\312' 0xCA
        " ## ",
        " ## ",
        "####",
        "####",
        "    ",
        "    ") &
      glyph( -- '\313' 0xCB
        "    ",
        "    ",
        "####",
        "####",
        " ## ",
        " ## ") &
      glyph( -- '\314' 0xCC
        " ## ",
        " ## ",
        " ###",
        " ###",
        " ## ",
        " ## ") &
      glyph( -- '\315' 0xCD
        "    ",
        "    ",
        "####",
        "####",
        "    ",
        "    ") &
      glyph( -- '\316' 0xCE
        " ## ",
        " ## ",
        "####",
        "####",
        " ## ",
        " ## ") &
      glyph( -- '\317' 0xCF
        "  # ",
        "  # ",
        "####",
        "####",
        "    ",
        "    ") &
      glyph( -- '\320' 0xD0
        " ## ",
        " ## ",
        "####",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\321' 0xD1
        "    ",
        "    ",
        "####",
        "####",
        "  # ",
        "  # ") &
      glyph( -- '\322' 0xD2
        "    ",
        "    ",
        "####",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\323' 0xD3
        " ## ",
        " ## ",
        " ###",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\324' 0xD4
        "  # ",
        "  # ",
        "  ##",
        "  ##",
        "    ",
        "    ") &
      glyph( -- '\325' 0xD5
        "    ",
        "    ",
        "  ##",
        "  ##",
        "  # ",
        "  # ") &
      glyph( -- '\326' 0xD6
        "    ",
        "    ",
        " ###",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\327' 0xD7
        " ## ",
        " ## ",
        "####",
        " ## ",
        " ## ",
        " ## ") &
      glyph( -- '\330' 0xD8
        "  # ",
        "  # ",
        "####",
        "####",
        "  # ",
        "  # ") &
      glyph( -- '\331' 0xD9
        "  # ",
        "  # ",
        "### ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\332' 0xDA
        "    ",
        "    ",
        "  ##",
        "  # ",
        "  # ",
        "  # ") &
      glyph( -- '\333' 0xDB
        "####",
        "####",
        "####",
        "####",
        "####",
        "####") &
      glyph( -- '\334' 0xDC
        "    ",
        "    ",
        "    ",
        "####",
        "####",
        "####") &
      glyph( -- '\335' 0xDD
        "##  ",
        "##  ",
        "##  ",
        "##  ",
        "##  ",
        "##  ") &
      glyph( -- '\336' 0xDE
        "  ##",
        "  ##",
        "  ##",
        "  ##",
        "  ##",
        "  ##") &
      glyph( -- '\337' 0xDF
        "####",
        "####",
        "####",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\340' 0xE0
        "    ",
        "    ",
        " # #",
        "# # ",
        " # #",
        "    ") &
      glyph( -- '\341' 0xE1
        " #  ",
        "# # ",
        "##  ",
        "# # ",
        "##  ",
        "#   ") &
      glyph( -- '\342' 0xE2
        "### ",
        "# # ",
        "#   ",
        "#   ",
        "#   ",
        "    ") &
      glyph( -- '\343' 0xE3
        "    ",
        "##  ",
        "# ##",
        "# # ",
        "# # ",
        "    ") &
      glyph( -- '\344' 0xE4
        "### ",
        "#   ",
        " #  ",
        "#   ",
        "### ",
        "    ") &
      glyph( -- '\345' 0xE5
        "    ",
        "    ",
        " ###",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- '\346' 0xE6
        "    ",
        "    ",
        "# # ",
        "# # ",
        "## #",
        "#   ") &
      glyph( -- '\347' 0xE7
        "    ",
        "##  ",
        " ###",
        " #  ",
        "  # ",
        "    ") &
      glyph( -- '\350' 0xE8
        " #  ",
        " #  ",
        "# # ",
        " #  ",
        "### ",
        "    ") &
      glyph( -- '\351' 0xE9
        " ## ",
        "# # ",
        "### ",
        "# # ",
        "##  ",
        "    ") &
      glyph( -- '\352' 0xEA
        " #  ",
        "# # ",
        "# # ",
        "# # ",
        "# ##",
        "    ") &
      glyph( -- '\353' 0xEB
        " ## ",
        "#   ",
        " #  ",
        "# # ",
        " ## ",
        "    ") &
      glyph( -- '\354' 0xEC
        "    ",
        "    ",
        " ## ",
        "### ",
        " ## ",
        "    ") &
      glyph( -- '\355' 0xED
        "    ",
        "    ",
        "   #",
        " ## ",
        " ## ",
        "#   ") &
      glyph( -- '\356' 0xEE
        " ###",
        "#   ",
        " ## ",
        "#   ",
        " ###",
        "    ") &
      glyph( -- '\357' 0xEF
        " ## ",
        "#  #",
        "#  #",
        "#  #",
        "#  #",
        "    ") &
      glyph( -- '\360' 0xF0
        "####",
        "    ",
        "####",
        "    ",
        "####",
        "    ") &
      glyph( -- '\361' 0xF1
        " #  ",
        "### ",
        " #  ",
        "    ",
        "### ",
        "    ") &
      glyph( -- '\362' 0xF2
        "#   ",
        " #  ",
        "### ",
        "    ",
        "### ",
        "    ") &
      glyph( -- '\363' 0xF3
        "  # ",
        " #  ",
        "### ",
        "    ",
        "### ",
        "    ") &
      glyph( -- '\364' 0xF4
        "  # ",
        " #  ",
        " #  ",
        " #  ",
        " #  ",
        " #  ") &
      glyph( -- '\365' 0xF5
        " #  ",
        " #  ",
        " #  ",
        " #  ",
        " #  ",
        "#   ") &
      glyph( -- '\366' 0xF6
        " #  ",
        "    ",
        "### ",
        "    ",
        " #  ",
        "    ") &
      glyph( -- '\367' 0xF7
        "##  ",
        "  ##",
        "    ",
        "##  ",
        "  ##",
        "    ") &
      glyph( -- '\370' 0xF8
        " ## ",
        "##  ",
        "    ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\371' 0xF9
        "    ",
        " #  ",
        "### ",
        " #  ",
        "    ",
        "    ") &
      glyph( -- '\372' 0xFA
        "    ",
        "    ",
        "  # ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\373' 0xFB
        "    ",
        "   #",
        "  # ",
        "# # ",
        " #  ",
        "    ") &
      glyph( -- '\374' 0xFC
        "##  ",
        "# # ",
        "# # ",
        "    ",
        "    ",
        "    ") &
      glyph( -- '\375' 0xFD
        "##  ",
        "  # ",
        "#   ",
        "### ",
        "    ",
        "    ") &
      glyph( -- '\376' 0xFE
        "    ",
        " ## ",
        " ## ",
        " ## ",
        " ## ",
        "    ") &
      glyph( -- '\377' 0xFF
        "    ",
        "    ",
        "    ",
        "    ",
        "    ",
        "    ")
      );

end package;
