library nsl_data;
use nsl_data.bytestream.all;

package neorv32_init is

  constant neorv32_bootrom_init : byte_string := from_hex(
    ""
    & "b7200000938000807390003097000000"
    & "9380c012739050307310403017210080"
    & "130101fe970100809381c17d13020000"
    & "93020000130300009303000013040000"
    & "93040000130800009308000013090000"
    & "93090000130a0000930a0000130b0000"
    & "930b0000130c0000930c0000130d0000"
    & "930d0000130e0000930e0000130f0000"
    & "930f0000971500009385454717060080"
    & "130646f7970600809386c6f6638ec500"
    & "635cd60003a705002320e60093854500"
    & "130646006ff0dffe17070080130787f4"
    & "938781806358f7002320070013074700"
    & "6ff05fff171400001304041897140000"
    & "93848417635a940083200400e7800000"
    & "130444006ff01fff1305000093050000"
    & "ef008007731040307310053417140000"
    & "130484149714000093840414635a9400"
    & "83200400e7800000130444006ff01fff"
    & "730050106ff0dfff7310043473242034"
    & "1354f401631604027324103413042400"
    & "731014347324a034137434001304d4ff"
    & "63080400732410341304240073101434"
    & "7324003473002030130101fd232c4101"
    & "370a008023220a00b707008023a00700"
    & "23261102232481022322910223202103"
    & "232e3101232a51012328610123267101"
    & "9307c06473905730ef00904a630e0500"
    & "13070000930600001306000093050000"
    & "13052000ef00d049ef00506d63040502"
    & "13052000130730009306000013060000"
    & "93050000ef00906cef00107913053000"
    & "ef009073ef00503c6308050013051000"
    & "93050000ef00503fb755000037f5ffff"
    & "13060000938505b013050550ef005052"
    & "ef00903e63080502b7f7ffff23a00740"
    & "23a20740032700e01357270023a4e740"
    & "23a60740930700087390473093078000"
    & "73a00730b715000037f5ffff93850539"
    & "13050550ef00d05c732530f1ef00c02c"
    & "b715000037f5ffff9385853c13050550"
    & "ef00105b032500e0ef00002bb7150000"
    & "37f5ffff9385053d13050550ef005059"
    & "73251030ef004029b715000037f5ffff"
    & "9385853d13050550ef009057732500fc"
    & "ef008027b715000037f5ffff9385053e"
    & "13050550ef00d055032580e013041000"
    & "37190000ef004025b715000037f5ffff"
    & "9385853e13050550ef009053034540e0"
    & "3315a4001375c5ffef000023b7150000"
    & "37f5ffff9385053f13050550ef005051"
    & "834750e03315f4001375c5ffef00c020"
    & "37f5ffff9305092f13050550ef00504f"
    & "ef00902c63080506b715000037f5ffff"
    & "9385853f13050550ef00904def00d02b"
    & "032400e0b7f9ffff9389095013143400"
    & "b304a40033b484003304b40013850900"
    & "ef0050386300050a13850900ef009048"
    & "630a050837f5ffff13050550ef009048"
    & "b715000037f5ffff9385454213050550"
    & "ef001048b7f4ffffb7190000ef004010"
    & "b71a000093840450130bf003930b3001"
    & "9389494893850a4313850400ef005045"
    & "13850400ef0090419305050013040500"
    & "13850400ef00903e9305092f13850400"
    & "ef0010436302640b1304b4f91374f40f"
    & "63e28b0a131424003304340183270400"
    & "67800700ef00501fe3ea85f46314b400"
    & "e36695f413051000ef00c05637f5ffff"
    & "9305092f13050550ef00903e13050000"
    & "ef000018b7c2ffff67800200ef004006"
    & "6ff05ff713050000ef00c0536ff09ff6"
    & "ef00c07a6ff01ff6130510006ff0dffe"
    & "83274a00e39407fcb715000093858543"
    & "37f5ffff13050550ef0090396ff09ff3"
    & "130510006ff0dffab715000093858544"
    & "6ff01ffeb7150000938585476ff05ffd"
    & "b715000037f5ffff9385452513050550"
    & "6f001036130101ff23248100b7150000"
    & "1304050037f5ffff9385452d13050550"
    & "23261100ef00d03393172400b7150000"
    & "b38787009385454e37f5ffffb385f500"
    & "13050550ef00d0319307800073b00730"
    & "ef009009630805001305100093050000"
    & "ef00900c6f000000130101fe23263101"
    & "9309050037f5ffff9305000313050550"
    & "232e1100232c8100232a910023282101"
    & "23244101ef00902737f5ffff93058007"
    & "1305055037190000b7f4ffffef001026"
    & "1304c0011309494d93840450130ac0ff"
    & "b3d7890093f7f700b307f90083c50700"
    & "138504001304c4ffef005023e31244ff"
    & "8320c101032481018324410103290101"
    & "8329c100032a81001301010267800000"
    & "130101ff232611002324810023229100"
    & "9307800073b007301304000063040500"
    & "370440e0b715000037f5ffff9385c52d"
    & "13050550ef00d02213050400eff0dff2"
    & "b715000037f5ffff9385c52e13050550"
    & "b7f4ffffef00d0209384045013850400"
    & "ef00101ce31c05fee7000400130101fb"
    & "23261104232451042322610423207104"
    & "232e8102232c9102232aa1022328b102"
    & "2326c1022324d1022322e1022320f102"
    & "232e0101232c1101232ac1012328d101"
    & "2326e1012324f101f3242034b7070080"
    & "938777006394f408ef00007263060500"
    & "13050000ef004072ef00007663000502"
    & "ef008076832700e093d727003385a700"
    & "b337f500b385b700ef00c0760324c103"
    & "8320c104832281040323410483230104"
    & "8324810303254103832501030326c102"
    & "8326810203274102832701020328c101"
    & "83288101032e4101832e0101032fc100"
    & "832f8100130101057300203093077000"
    & "639cf400b707008083a7070063860700"
    & "13051000eff01fda7324103437f5ffff"
    & "13050550ef00007c63020506b7150000"
    & "37f5ffff9385452f13050550ef00500d"
    & "13850400eff05fdd37f5ffff93050002"
    & "13050550ef00900613050400eff0dfdb"
    & "37f5ffff9305000213050550ef001005"
    & "73253034eff05fdab715000037f5ffff"
    & "9385052f13050550ef00900813044400"
    & "731014346ff09ff1130101ff13050000"
    & "23261100ef00006f1305b00aef000072"
    & "8320c100130101016f000070130101ff"
    & "1305000023261100ef00c06c13056000"
    & "ef00c06f8320c100130101016f00c06d"
    & "130101ff1305000023261100ef00806a"
    & "13054000ef00806d8320c10013010101"
    & "6f00806b130101fe13050000232e1100"
    & "ef00406813055000ef00406b13050000"
    & "ef00c06a2326a100ef0000698320c101"
    & "0325c1001301010267800000130101ff"
    & "23261100eff05ff5eff05ff7eff09ffb"
    & "937725001305f0ff638a0700eff05ff8"
    & "eff05ffa1315e5011355f5418320c100"
    & "1301010167800000130101ff23248100"
    & "13040500135505011375f50f23261100"
    & "ef00c063135584001375f50fef000063"
    & "1375f40f032481008320c10013010101"
    & "6f00c061130101fe232c810013040500"
    & "13050000232e1100ef00c05c13053000"
    & "ef00c05f13050400eff01ffa13050000"
    & "ef00c05e2326a100ef00005d8320c101"
    & "032481010325c1001301010267800000"
    & "130101fd232e3101b7f9ffff23248102"
    & "2322910223202103232c410123261102"
    & "93040500138905001304000093890950"
    & "130a40006392040413850900ef00006a"
    & "9307c100b38787002380a70013041400"
    & "e31244ff8320c102032481020325c100"
    & "83244102032901028329c101032a8101"
    & "130101036780000033058900eff09ff3"
    & "6ff01ffc130101fd2328610193071000"
    & "370b0080232481022326110223229102"
    & "23202103232e3101232c4101232a5101"
    & "232671012320fb0013040500631c0502"
    & "b715000037f5ffff9385053013050550"
    & "ef000064b705400013050400eff05ff2"
    & "b7d788479387e7af630ef50413050000"
    & "6f004004b715000037f5ffff93850532"
    & "13050550ef00c06037054000eff0dfb0"
    & "b715000037f5ffff9385c53213050550"
    & "ef00005f832780e01397d70063460700"
    & "13053000eff01fa8eff05fe0e30c05f8"
    & "6ff01fffb70540009385450013050400"
    & "eff01febb70540009309050093858500"
    & "13050400eff0dfe9b70a4000130a0500"
    & "93fbc9ff1309000093040000938aca00"
    & "b3055901631e7905b384440113052000"
    & "e39204fab715000037f5ffff93854533"
    & "13050550ef00c0568320c10203248102"
    & "b707008023a2370123200b0083244102"
    & "032901028329c101032a8101832a4101"
    & "032b0101832bc1001301010367800000"
    & "13050400eff0dfe12320a900b384a400"
    & "130949006ff0dff8130101ff23261100"
    & "23248100232291001384050093040500"
    & "eff0dfca13050000ef00c03713052000"
    & "ef00c03a13850400eff01fd513050400"
    & "ef00c039ef004038eff0dfcc13751500"
    & "e31c05fe8320c1000324810083244100"
    & "1301010167800000130101fe232c8100"
    & "232a910023282101232e110093040500"
    & "2326b10013040000130940009307c100"
    & "b387870083c507003385840013041400"
    & "eff09ff6e31424ff8320c10103248101"
    & "83244101032901011301010267800000"
    & "130101ff232611002324810013040500"
    & "eff0dfbf13050000ef00c02c1305800d"
    & "ef00c02f13050400eff01fcaef00c02d"
    & "eff05fc213751500e31c05fe8320c100"
    & "032481001301010167800000130101fe"
    & "b7070080232c810003a44700232e1100"
    & "232a9100232821012326310123244101"
    & "631a0402b71500009385853303248101"
    & "8320c10183244101032901018329c100"
    & "032a810037f5ffff1305055013010102"
    & "6f00003cb715000037f5ffff93854535"
    & "13050550ef00c03a13050400eff0df8a"
    & "b715000037f5ffff9385c53513050550"
    & "ef00003937054000eff01f89b7150000"
    & "37f5ffff9385453713050550ef004037"
    & "37f5ffff13050550ef00403393050500"
    & "9304050037f5ffff13050550ef000030"
    & "93079007639af40aeff05fb763060500"
    & "13053000eff00ffeb715000037f5ffff"
    & "9385053813050550ef00803293540401"
    & "37094000370a01009309f0ff13050900"
    & "9384f4ffeff0dfea33094901e39834ff"
    & "b709400093040000130900009389c900"
    & "9387040083a507003385340193844400"
    & "3309b900eff05fe2e3e484feb7d58847"
    & "9385e5af37054000eff01fe137054000"
    & "9305040013054500eff01fe037054000"
    & "b305204113058500eff01fdfb7150000"
    & "938545336ff09feb8320c10103248101"
    & "83244101032901018329c100032a8100"
    & "1301010267800000032580e01355f500"
    & "1375150067800000930710001307f001"
    & "b397a700634aa700032780c0b347f700"
    & "2324f0c0678000000327c0c0b347f700"
    & "2326f0c067800000930700c023a4a700"
    & "23a6b70067800000032580e013550501"
    & "1375150067800000b7f7ffff93870740"
    & "83a5470003a5070003a74700e39ae5fe"
    & "67800000b7f7ffff1307f0ff23a4e740"
    & "23a6b74023a4a7401300000067800000"
    & "032580e0135525011375150067800000"
    & "b70770003377f70013161600b7470000"
    & "137626009395a500938707c03366e600"
    & "b3f5f500131575003366b60013750538"
    & "939626003366a60093f6460013080080"
    & "3366d60023200800136616002320c800"
    & "678000009306008003a7060093173500"
    & "93f78703137777f8b3e7e70093e70704"
    & "23a0f600678000001307008083270700"
    & "93f7f7fb2320f700678000002322a080"
    & "83270080e3ce07fe032540801375f50f"
    & "6780000037f7ffff1307075093070500"
    & "631ae500032580e01355150113751500"
    & "6780000037f7ffff1307076013050000"
    & "e398e7fe032580e0135595016ff01ffe"
    & "130101ff232481002322910023261100"
    & "2320050093040500032500e093951500"
    & "13040600ef004023130700009306e03f"
    & "63e6a6049307f5ffb7060100938606fc"
    & "93976700b3f7d700b706c0073374d400"
    & "13173700b3e78700137787018320c100"
    & "03248100b3e7e70093e7170023a0f400"
    & "8324410013010101678000009307e7ff"
    & "93f7d7ff639807001355350013071700"
    & "6ff01ffa135515006ff05fff83270500"
    & "1397a700e34c07fe2322b50067800000"
    & "032505001355f5016780000083270500"
    & "1397f700e35c07fe032545001375f50f"
    & "67800000032505001355050113751500"
    & "67800000032545001375f50f67800000"
    & "130101fe232c8100232a910023263101"
    & "232e1100232821019304050013840500"
    & "9309a000034904001304140063100902"
    & "8320c101032481018324410103290101"
    & "8329c100130101026780000063183901"
    & "9305d00013850400eff05ff593050900"
    & "13850400eff09ff46ff0dffb032580e0"
    & "1355d501137515006780000093958501"
    & "3708000fb3f505011317d70093965600"
    & "b7f7ffffb3e5e50093f6060213164600"
    & "b3e5d500137606011315150023a007f0"
    & "b3e5c5001375e50023a407f0b3e5a500"
    & "23a607f093e5152023a0b7f023a407f0"
    & "938707f023a6070003a7070093161700"
    & "e3cc06fe03a70700b70620003367d700"
    & "23a0e700678000009307f5ff13073000"
    & "6360f70437f7ffff832607f037e6ffff"
    & "1306f67fb3f6c6009397b700b3e7d700"
    & "1305550093f7f7c3131565003365f500"
    & "136505402320a7f01305000067800000"
    & "1305f0ff67800000b7f7ffff03a707f0"
    & "b70680003367d70023a0e7f067800000"
    & "6340050663c605061386050093050500"
    & "1305f0ff630c060293061000637ab600"
    & "6358c0001316160093961600e36ab6fe"
    & "1305000063e6c500b385c5403365d500"
    & "93d6160013561600e39606fe67800000"
    & "93820000eff05ffb1385050067800200"
    & "3305a0406348b000b305b0406ff0dff9"
    & "b305b04093820000eff01ff93305a040"
    & "678002009382000063ca0500634c0500"
    & "eff09ff71385050067800200b305b040"
    & "e35805fe3305a040eff01ff63305b040"
    & "67800200417661696c61626c6520434d"
    & "44733a0a20683a2048656c700a20723a"
    & "20526573746172740a20753a2055706c"
    & "6f61640a20733a2053746f726520746f"
    & "20666c6173680a206c3a204c6f616420"
    & "66726f6d20666c6173680a20783a2042"
    & "6f6f742066726f6d20666c6173682028"
    & "584950290a20653a2045786563757465"
    & "00000000070a4552525f0000426f6f74"
    & "696e672066726f6d200000002e2e2e0a"
    & "0a0000000a4552525f45584320000000"
    & "4177616974696e67206e656f72763332"
    & "5f6578652e62696e2e2e2e2000000000"
    & "4c6f6164696e672028400000292e2e2e"
    & "0a0000004f4b00004e6f206578656375"
    & "7461626c6520617661696c61626c652e"
    & "00000000577269746520000020627974"
    & "657320746f2053504920666c61736820"
    & "402000003f2028792f6e292000000000"
    & "0a466c617368696e672e2e2e20000000"
    & "0a0a0a3c3c204e454f5256333220426f"
    & "6f746c6f61646572203e3e0a0a424c44"
    & "563a204a616e20323120323032340a48"
    & "57563a20200000000a434c4b3a202000"
    & "0a4d4953413a20000a584953413a2000"
    & "0a534f433a2020000a494d454d3a2000"
    & "0a444d454d3a20000a4175746f626f6f"
    & "7420696e2038732e2050726573732061"
    & "6e79206b657920746f2061626f72742e"
    & "0a00000041626f727465642e0a0a0000"
    & "0a434d443a3e20004e6f206578656375"
    & "7461626c652e00006279205374657068"
    & "616e204e6f6c74696e670a6769746875"
    & "622e636f6d2f73746e6f6c74696e672f"
    & "6e656f7276333200496e76616c696420"
    & "434d440090040000c4040000c4040000"
    & "6c040000c4040000c4040000c4040000"
    & "88040000c4040000c4040000c4040000"
    & "c4040000c40400006404000080040000"
    & "c404000074040000c4040000c4040000"
    & "b0040000303132333435363738396162"
    & "63646566455845000053495a45004348"
    & "4b5300464c534800"
    );
  constant neorv32_imem_init : byte_string := null_byte_string;

end package neorv32_init;
