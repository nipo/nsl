library ieee;
use ieee.std_logic_1164.all;

library nsl;

entity framed_spi_controller is
  generic(
    slave_count   : natural range 1 to 63 := 1
    );
  port(
    clock : in std_logic;
    resetn : in std_logic;

    framed_cmd_data : in std_logic_vector(7 downto 0);
    framed_cmd_last : in std_logic;
    framed_cmd_valid : in std_logic;
    framed_cmd_ready : out std_logic;
    framed_rsp_data : out std_logic_vector(7 downto 0);
    framed_rsp_last : out std_logic;
    framed_rsp_valid : out std_logic;
    framed_rsp_ready : in std_logic;

    spi_cs_n : out std_logic_vector(0 to slave_count-1);
    spi_sck : out std_logic;
    spi_mosi : out std_logic;
    spi_miso : in std_logic
    );
end entity;

architecture rtl of framed_spi_controller is

  -- attributes for ports should be in entity block, and case is supposed to be
  -- non-sensitive, but Xilinx tools only take upper-cased names attributes,
  -- and only if they are inside the architecture block... Go figure.
  attribute X_INTERFACE_INFO : string;
  attribute X_INTERFACE_PARAMETER : string;

  attribute X_INTERFACE_PARAMETER of clock : signal is "ASSOCIATED_BUSIF framed, ASSOCIATED_RESET resetn";
  attribute X_INTERFACE_PARAMETER of resetn : signal is "POLARITY ACTIVE_LOW";

  attribute X_INTERFACE_INFO of framed_cmd_ready : signal is "nsl:interface:framed:1.0 framed req_ready";
  attribute X_INTERFACE_INFO of framed_cmd_valid : signal is "nsl:interface:framed:1.0 framed req_valid";
  attribute X_INTERFACE_INFO of framed_cmd_last  : signal is "nsl:interface:framed:1.0 framed req_last";
  attribute X_INTERFACE_INFO of framed_cmd_data  : signal is "nsl:interface:framed:1.0 framed req_data";
  attribute X_INTERFACE_INFO of framed_rsp_ready : signal is "nsl:interface:framed:1.0 framed rsp_ready";
  attribute X_INTERFACE_INFO of framed_rsp_valid : signal is "nsl:interface:framed:1.0 framed rsp_valid";
  attribute X_INTERFACE_INFO of framed_rsp_last  : signal is "nsl:interface:framed:1.0 framed rsp_last";
  attribute X_INTERFACE_INFO of framed_rsp_data  : signal is "nsl:interface:framed:1.0 framed rsp_data";

  attribute X_INTERFACE_INFO of spi_cs_n : signal is "nsl:interface:spi:1.0 spi cs_n";
  attribute X_INTERFACE_INFO of spi_sck  : signal is "nsl:interface:spi:1.0 spi sck";
  attribute X_INTERFACE_INFO of spi_miso : signal is "nsl:interface:spi:1.0 spi miso";
  attribute X_INTERFACE_INFO of spi_mosi : signal is "nsl:interface:spi:1.0 spi mosi";

  signal rsp_data : std_ulogic_vector(7 downto 0);
  
begin

  controller: nsl.spi.spi_master
    generic map(
      slave_count => slave_count
      )
    port map(
      p_resetn => resetn,
      p_clk => clock,

      p_cmd_val.valid => framed_cmd_valid,
      p_cmd_val.data => std_ulogic_vector(framed_cmd_data),
      p_cmd_val.last => framed_cmd_last,
      p_cmd_ack.ready => framed_cmd_ready,
      p_rsp_val.valid => framed_rsp_valid,
      p_rsp_val.data => rsp_data,
      p_rsp_val.last => framed_rsp_last,
      p_rsp_ack.ready => framed_rsp_ready,

      p_sck => spi_sck,
      std_logic_vector(p_csn) => spi_cs_n,
      p_mosi => spi_mosi,
      p_miso => spi_miso
      );

  framed_rsp_data <= std_logic_vector(rsp_data);
  
end;
