library ieee;
use ieee.std_logic_1164.all;

package pmod is
  
  subtype pmod_io_t is std_logic_vector(0 to 7);

end package pmod;
