package control is

  procedure terminate(retval : integer);
  
end package control;
