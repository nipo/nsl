library nsl_data;
use nsl_data.bytestream.all;



-- Extracted from:
-- 
-- - main.elf
--   ElfProgram:
--    + device: RISC-V
--    + entry: 0xffffc000 (4294950912)
--    - <0xffffc000:0xffffcda0 (3488 bytes) '.text .rodata'>
--    - <0xffffcd98:0xffffcda0 (8 bytes) '.bss'>

package neorv32_bootrom is


  constant init : byte_string := from_hex(""
    & "b72000009380008073900030970000009380c012739050307310403017410080"
    & "1301011e974100809381c17d1302000093020000130300009303000013040000"
    & "9304000013080000930800001309000093090000130a0000930a0000130b0000"
    & "930b0000130c0000930c0000130d0000930d0000130e0000930e0000130f0000"
    & "930f000097150000938545d117460080130646f7974600809386c6f6638ec500"
    & "635cd60003a705002320e60093854500130646006ff0dffe17470080130787f4"
    & "938781806358f70023200700130747006ff05fff17140000130444b397140000"
    & "9384c4b2635a940083200400e7800000130444006ff01fff1305000093050000"
    & "ef0080077310403073100534171400001304c4af97140000938444af635a9400"
    & "83200400e7800000130444006ff01fff730050106ff0dfff7310043473242034"
    & "1354f401631604027324103413042400731014347324a034137434001304d4ff"
    & "630804007324103413042400731014347324003473002030130101fb23202105"
    & "37090080232e310323220900b7090080b7c7ffff232611042324810423229104"
    & "232c4103232a5103232861032326710323248103232291032320a103232eb101"
    & "23a009009387476573905730ef00500963040502130520001307300093060000"
    & "1306000093050000ef009008ef00101513053000ef00900fef00406463080500"
    & "1305100093050000ef004067b7c5010037f5ffff130600009385052013050550"
    & "ef00006f37f5ffff13050550ef000078ef00c06563080502b7f7ffff23a00740"
    & "23a20740032700e01357270023a4e74023a60740930700087390473093078000"
    & "73a00730b7d5ffff37f5ffff938585c313050550ef000078732530f1ef000028"
    & "b7d5ffff37f5ffff938505c713050550ef004076032500e0ef004026b7d5ffff"
    & "37f5ffff938585c713050550ef00807473251030ef008024b7d5ffff37f5ffff"
    & "938505c813050550ef00c072732500fcef00c022b7d5ffff37f5ffff938585c8"
    & "13050550ef000071032580e01304100037daffffef008020b7d5ffff37f5ffff"
    & "938505c913050550ef00c06e034540e0b7daffffb7f4ffff3315a4001375c5ff"
    & "ef00c01db7d5ffff37f5ffff938585c913050550ef00006c834750e0b7dbffff"
    & "938404503315f4001375c5ffef00001b37f5ffff9305cac113050550ef008069"
    & "b7d5ffff37f5ffff938505ca13050550ef00406837f5ffff93854aca13050550"
    & "ef004067130b8006130c5007930c8007130df003930d50069385cbcf13850400"
    & "ef00406513850400ef004063930505001304050013850400ef0040609305cac1"
    & "13850400ef000063630a6403636c8b006300a413630cb40fb7d5ffff938585d6"
    & "6f000002630684036300941193072007e314f4feb7c2ffff6780020093854aca"
    & "37f5ffff13050550ef00c05e6ff0dff8b7d5ffff37f5ffff93071000938545d0"
    & "1305055023a0f900ef00c05cef008016b7d788479387e7af6306f50013050000"
    & "ef00001bef00001513040500ef00801493070500135624001307000093060000"
    & "631ac700b387d70063820704130520006ff01ffd2326c1002324e1002322d100"
    & "2320f100ef00001103278100832641000326c1009315270083270100b386a600"
    & "23a0a500130717006ff09ffbb7d5ffff37f5ffff938545d213050550ef008053"
    & "2322890023a009006ff01fed8327490063980700b7d5ffff938585d26ff05ff2"
    & "13050000ef00c02e130510006ff09fffb7d5ffff938585d36ff09ff0130101fe"
    & "232631019309050037f5ffff9305000313050550232e1100232c8100232a9100"
    & "2328210123244101ef00404937f5ffff930580071305055037d9ffffb7f4ffff"
    & "ef00c0471304c001130949d793840450130ac0ffb3d7890093f7f700b307f900"
    & "83c50700138504001304c4ffef000045e31244ff8320c1010324810183244101"
    & "032901018329c100032a81001301010267800000130101fe232a9100b7f4ffff"
    & "232c810023282101232e110013040000938404501309400013850400ef000042"
    & "9307c100b38787002380a70013041400e31424ff8320c101032481010325c100"
    & "83244101032901011301010267800000130101ff23248100b7d5ffff13040500"
    & "37f5ffff938585c01305055023261100ef00403e93172400b7d5ffffb3878700"
    & "938545d837f5ffffb385f50013050550ef00403c9307800073b00730ef000020"
    & "630805001305100093050000ef0000236f000000130101fb2326110423245104"
    & "2322610423207104232e8102232c9102232aa1022328b1022326c1022324d102"
    & "2322e1022320f102232e0101232c1101232ac1012328d1012326e1012324f101"
    & "f3242034b7070080938777006394f408ef00c0186306050013050000ef000019"
    & "ef00c01c63000502ef00401d832700e093d727003385a700b337f500b385b700"
    & "ef00801d0324c1038320c1048322810403234104832301048324810303254103"
    & "832501030326c1028326810203274102832701020328c10183288101032e4101"
    & "832e0101032fc100832f8100130101057300203093077000639cf400b7070080"
    & "83a707006386070013051000eff05fea7324103437f5ffff13050550ef008017"
    & "63020506b7d5ffff37f5ffff938505c113050550ef00002813850400eff01fd8"
    & "37f5ffff9305000213050550ef00002313050400eff09fd637f5ffff93050002"
    & "13050550ef00802173253034eff01fd5b7d5ffff37f5ffff9385c5c113050550"
    & "ef00402313044400731014346ff09ff1130101ff232611002324810023229100"
    & "9307800073b007301304000063040500370440e0b7d5ffff37f5ffff938505c2"
    & "13050550ef00001f13050400eff01fcfb7d5ffff37f5ffff938505c313050550"
    & "b7f4ffffef00001d9384045013850400ef00001ae31c05fee7000400032580e0"
    & "1355f5001375150067800000930710001307f001b397a700634aa700032780c0"
    & "b347f7002324f0c0678000000327c0c0b347f7002326f0c067800000930700c0"
    & "23a4a70023a6b70067800000032580e0135505011375150067800000b7f7ffff"
    & "9387074083a5470003a5070003a74700e39ae5fe67800000b7f7ffff1307f0ff"
    & "23a4e74023a6b74023a4a740130000006780000037f7ffff1307075093070500"
    & "631ae500032580e013551501137515006780000037f7ffff1307076013050000"
    & "e398e7fe032580e0135595016ff01ffe130101ff232481002322910023261100"
    & "2320050093040500032500e09395150013040600ef008022130700009306e03f"
    & "63e6a6049307f5ffb7060100938606fc93976700b3f7d700b706c0073374d400"
    & "13173700b3e78700137787018320c10003248100b3e7e70093e7170023a0f400"
    & "8324410013010101678000009307e7ff93f7d7ff639807001355350013071700"
    & "6ff01ffa135515006ff05fff8327050093e747002320f5006780000083270500"
    & "1397a700e34c07fe2322b50067800000032505001355f5016780000083270500"
    & "1397f700e35c07fe032545001375f50f67800000130101fe232c8100232a9100"
    & "23263101232e11002328210193040500138405009309a0000349040013041400"
    & "631009028320c1010324810183244101032901018329c1001301010267800000"
    & "631839019305d00013850400eff01ff79305090013850400eff05ff66ff0dffb"
    & "032580e01355d5011375150067800000939585013708000fb3f505011317d700"
    & "93965600b7f7ffffb3e5e50093f6060213164600b3e5d5001376060113151500"
    & "23a007f0b3e5c5001375e50023a407f0b3e5a50023a607f093e5152023a0b7f0"
    & "23a407f0938707f023a6070003a7070093161700e3cc06fe03a70700b7062000"
    & "3367d70023a0e700678000009307f5ff130730006360f70437f7ffff832607f0"
    & "37e6ffff1306f67fb3f6c6009397b700b3e7d7001305550093f7f7c313156500"
    & "3365f500136505402320a7f013050000678000001305f0ff67800000b7f7ffff"
    & "03a707f0b70680003367d70023a0e7f0678000006340050663c6050613860500"
    & "930505001305f0ff630c060293061000637ab6006358c0001316160093961600"
    & "e36ab6fe1305000063e6c500b385c5403365d50093d6160013561600e39606fe"
    & "6780000093820000eff05ffb13850500678002003305a0406348b000b305b040"
    & "6ff0dff9b305b04093820000eff01ff93305a040678002009382000063ca0500"
    & "634c0500eff09ff71385050067800200b305b040e35805fe3305a040eff01ff6"
    & "3305b04067800200070a4552525f00000a4552525f455843200000000a000000"
    & "426f6f74696e672066726f6d200000002e2e2e0a0a0000000a0a0a3c3c204e45"
    & "4f5256333220426f6f746c6f61646572203e3e0a0a424c44563a204a616e2032"
    & "3420323032340a4857563a20200000000a434c4b3a2020000a4d4953413a2000"
    & "0a584953413a20000a534f433a2020000a494d454d3a20000a444d454d3a2000"
    & "0a0a0000417661696c61626c6520434d44733a0a20683a2048656c700a20723a"
    & "20526573746172740a20753a2055706c6f61640a20783a20426f6f742066726f"
    & "6d20666c6173682028584950290a20653a20457865637574650000000a434d44"
    & "3a3e20004177616974696e67206e656f727633325f6578652e62696e2e2e2e20"
    & "000000004f4b00004e6f2065786563757461626c652e00006279205374657068"
    & "616e204e6f6c74696e670a6769746875622e636f6d2f73746e6f6c74696e672f"
    & "6e656f7276333200496e76616c696420434d4400303132333435363738396162"
    & "63646566455845000053495a450043484b5300464c5348000000000000000000"
  );

end package neorv32_bootrom;
