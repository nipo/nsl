library ieee;
use ieee.std_logic_1164.all;

package types is
  
  subtype nsl_id is std_ulogic_vector(3 downto 0);
  
end package types;
