library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library nsl_data, nsl_amba, nsl_math, nsl_logic;
use nsl_data.bytestream.all;
use nsl_amba.axi4_stream.all;
use nsl_amba.random_pkt_checker.all;
use nsl_data.crc.all;
use nsl_data.prbs.all;
use nsl_logic.bool.all;

entity random_pkt_validator is
  generic (
    mtu_c: integer := 1500;
    config_c: config_t;
    data_prbs_init: prbs_state := x"deadbee"&"111";
    data_prbs_poly: prbs_state := prbs31;
    header_crc_params_c: crc_params_t
    );
  port (
    clock_i : in std_ulogic;
    reset_n_i : in std_ulogic;
    --
    in_i : in master_t;
    in_o : out slave_t;
    --
    out_o : out master_t;
    out_i : in slave_t
    );
end entity;

architecture beh of random_pkt_validator is

    constant header_config_c : buffer_config_t := buffer_config(config_c, HEADER_SIZE);
    constant max_nbr_data_cycle_l2 : integer := nsl_math.arith.log2(mtu_c/config_c.data_width);
    constant data_width_l2 : integer := nsl_math.arith.log2(config_c.data_width);
    constant stats_buf_config : buffer_config_t := buffer_config(config_c, STATS_SIZE);
    constant header_size_m1 : integer := HEADER_SIZE - 1;
    constant header_size_m_data_width : integer := HEADER_SIZE - config_c.data_width;
    constant stats_reset : stats_t := (
                                        stats_seqnum        => to_unsigned(0, 16),
                                        stats_pkt_size      => to_unsigned(0, 16),
                                        stats_header_valid  => true,
                                        stats_payload_valid => true,
                                        stats_index_data_ko => to_unsigned(0, 16)
                                    );

    function compare_with_keep(
        expected : byte_string;
        actual   : byte_string;
        keep     : std_ulogic_vector
      ) return boolean is
      begin
        for i in expected'range loop
          if keep(i) = '1' then
            if expected(i) /= actual(i) then
              return false;
            end if;
          end if;
        end loop;
        return true;
      end function;
      
    type state_t is (
        ST_RESET,
        ST_HEADER_DEC,
        ST_REALIGN_BUF,
        ST_HEADER_STATS,
        ST_DATA,
        ST_SEND_STATS_NO_EOP,
        ST_SEND_STATS_EOP,        
        ST_RESET_STATS
        );

    type txer_stats_t is (
        TXER_IDLE,
        TXER_SEND_STATS
        ); 

    type regs_t is
        record
            state : state_t;
            txer : txer_stats_t;
            state_pkt_gen :  prbs_state(30 downto 0);
            rx_bytes : unsigned(15 downto 0);
            header_buf : buffer_t;
            stats : stats_t;
            stats_buf : buffer_t;
            header : header_t;
            header_index_ko : integer range 0 to HEADER_SIZE - 1;
            seq_num : unsigned(15 downto 0);
            realign_cnt : integer range 0 to header_config_c.data_width;
            -- 
            header_valid_vector_debug : std_ulogic_vector(3 downto 0);
            payload_ref_debug : byte_string(0 to config_c.data_width -1);
            header_byte_debug : byte_string(0 to HEADER_SIZE-1);
            header_ref_byte_debug : byte_string(0 to HEADER_SIZE-1);
        end record;

    signal r, rin: regs_t;

begin
    regs: process(reset_n_i, clock_i) is
    begin
      if rising_edge(clock_i) then
        r <= rin;
      end if;
      if reset_n_i = '0' then
        r.state <= ST_RESET;
        r.txer <= TXER_IDLE;
        r.state_pkt_gen <= data_prbs_init;
        r.header_buf <= reset(header_config_c);
        r.stats_buf <= reset(stats_buf_config);
        r.rx_bytes <= (others => '0');
        r.seq_num <= (others => '0');
        r.stats.stats_seqnum <= (others => '0');
        r.stats.stats_pkt_size <= (others => '0');
        r.stats.stats_header_valid <= true;
        r.stats.stats_payload_valid <= true;
        r.header_index_ko <= 0;
        r.stats.stats_index_data_ko <= (others => '0');
        r.realign_cnt <= 0;
      end if;
    end process;

    rx_process: process(r, in_i, out_i, rin, clock_i)
        variable header : header_t;
        variable next_header_byte_string,header_byte_string : byte_string(0 to HEADER_SIZE-1);
        variable header_valid_v : boolean;
        variable payload_byte_ref_v : byte_string(0 to config_c.data_width -1);
        variable header_byte_ref_v, rx_header_v : byte_string(0 to HEADER_SIZE-1);
        variable send_stats_trigger_v : boolean;
    begin
        rin <= r;

        header := header_unpack(bytes(header_config_c,r.header_buf), to_integer(r.rx_bytes));
        rx_header_v := bytes(header_config_c,r.header_buf);

        next_header_byte_string := bytes(header_config_c,shift(header_config_c, r.header_buf, in_i));
        header_byte_string := bytes(header_config_c,r.header_buf);

        header_byte_ref_v := ref_header(r.rx_bytes,
                                        header,
                                        r.seq_num,
                                        header_crc_params_c);

        header_valid_v := is_header_valid(r.rx_bytes,
                                          header,
                                          r.seq_num,
                                          header_crc_params_c);

        payload_byte_ref_v := prbs_byte_string(r.state_pkt_gen, 
                                           data_prbs_poly,
                                           config_c.data_width);

        send_stats_trigger_v := false;

        case r.state is

            when ST_RESET =>
                rin.state <= ST_HEADER_DEC;

            when ST_HEADER_DEC =>
                if is_valid(config_c, in_i) then
                    rin.header_buf <= shift(header_config_c, r.header_buf, in_i);
                    rin.rx_bytes <= r.rx_bytes + count_valid_bytes(keep(config_c, in_i));
                    rin.stats.stats_payload_valid <= true;
                    if is_last(header_config_c, r.header_buf) or is_last(config_c, in_i) then
                        rin.seq_num <= r.seq_num + 1;
                        if should_align(header_config_c, r.header_buf,in_i) then
                            rin.realign_cnt <= header_config_c.beat_count - beat_count(header_config_c, shift(header_config_c, r.header_buf, in_i));
                            rin.state <= ST_REALIGN_BUF;
                        else
                            rin.state <= ST_HEADER_STATS;
                        end if;
                    end if;
                end if;

                when ST_REALIGN_BUF => 
                    if r.realign_cnt /= 0 then
                        rin.header_buf <= realign(header_config_c, r.header_buf);
                        rin.realign_cnt <= r.realign_cnt - 1;
                    else
                        rin.state <= ST_HEADER_STATS;
                    end if;

                when ST_HEADER_STATS =>
                    if header.pkt_size <= HEADER_SIZE then
                        rin.state <= ST_RESET_STATS;
                    else
                        rin.state <= ST_DATA;
                    end if;
                    --
                    for i in 0 to to_integer(r.rx_bytes) - 1 loop
                        if header_byte_ref_v(i) /= rx_header_v(i) then
                            rin.stats.stats_header_valid <= false;
                            rin.stats.stats_index_data_ko <= to_unsigned(i,r.stats.stats_index_data_ko'length);
                            rin.header_index_ko <= i;              
                            if header.pkt_size <= HEADER_SIZE then
                                rin.state <= ST_SEND_STATS_EOP;
                            else
                                rin.state <= ST_SEND_STATS_NO_EOP;
                            end if;
                            --
                            exit;
                        end if;
                    end loop;
                    rin.header <= header;
                    rin.stats.stats_seqnum <= header.seq_num;
                    rin.stats.stats_pkt_size <= header.pkt_size;
                    --
                    rin.header_byte_debug <= rx_header_v;
                    rin.header_ref_byte_debug <= header_byte_ref_v;
                    rin.header_valid_vector_debug <= is_header_valid_vector(r.rx_bytes,
                                                                           header,
                                                                           r.seq_num,
                                                                           header_crc_params_c);

                when ST_DATA => 
                    if is_valid(config_c, in_i) then
                        rin.rx_bytes <= r.rx_bytes + count_valid_bytes(keep(config_c, in_i));
                        rin.payload_ref_debug <= payload_byte_ref_v;
                        rin.state_pkt_gen <= prbs_forward(r.state_pkt_gen, 
                                                        data_prbs_poly,
                                                        count_valid_bytes(keep(config_c, in_i)) * 8);
                        --
                        for i in payload_byte_ref_v'range loop
                            if keep(config_c, in_i)(i) = '1' then
                                if payload_byte_ref_v(i) /= bytes(config_c, in_i)(i) then
                                    rin.stats.stats_payload_valid <= false;
                                    rin.stats.stats_index_data_ko <= r.rx_bytes + i;   
                                    send_stats_trigger_v := true;                           
                                  end if;
                            end if;
                          end loop;
                        --
                        if is_last(config_c, in_i) then
                            rin.state <= ST_RESET_STATS;
                            --
                            -- This distinction is necessary in the case of an inserted error in the 
                            -- packet size. Since we use the received packet size field to generate 
                            -- a reference header, an error inserted in this field will be detected 
                            -- in the random data and not directly in the size field.
                            --
                            if not (r.header_index_ko = 4 or r.header_index_ko = 5) then -- Test if error is in rand filed so in size field
                                if r.rx_bytes + count_valid_bytes(keep(config_c, in_i)) /= header.pkt_size then
                                    rin.stats.stats_payload_valid <= false;
                                    send_stats_trigger_v := true;                           
                                end if;
                            end if;
                        end if;
                        --
                        if send_stats_trigger_v then
                            rin.state <= ST_SEND_STATS_NO_EOP;
                            if is_last(config_c, in_i) then
                                rin.state <= ST_SEND_STATS_EOP;
                            end if;
                        end if;
                    end if;

                when ST_RESET_STATS => 
                    if r.txer = TXER_IDLE then
                        rin.stats_buf <= reset(stats_buf_config);
                        rin.header_buf <= reset(header_config_c);
                        rin.rx_bytes <= (others => '0');
                        rin.stats <= stats_reset;
                        rin.state <= ST_HEADER_DEC;
                    end if;

                when ST_SEND_STATS_NO_EOP => 
                    if r.txer = TXER_IDLE then
                        rin.stats_buf <= reset(stats_buf_config,stats_pack(r.stats));
                        if r.txer = TXER_IDLE then
                            rin.stats.stats_payload_valid <= true;
                            rin.state <= ST_DATA;
                        end if;
                    end if;         
     
                when ST_SEND_STATS_EOP => 
                    if r.txer = TXER_IDLE then
                        rin.stats_buf <= reset(stats_buf_config,stats_pack(r.stats));
                        rin.header_buf <= reset(header_config_c);
                        rin.rx_bytes <= (others => '0');
                        rin.stats <= stats_reset;
                        rin.state <= ST_HEADER_DEC;
                    end if;               

            when others => 
        end case;

        case r.txer is 
            when TXER_IDLE =>
                if r.state = ST_SEND_STATS_EOP or r.state = ST_SEND_STATS_NO_EOP then
                    rin.txer <= TXER_SEND_STATS;
                end if;

            when TXER_SEND_STATS =>
                if is_ready(config_c, out_i) then
                    rin.stats_buf <= shift(stats_buf_config, r.stats_buf);
                    if is_last(stats_buf_config, r.stats_buf) then
                        rin.txer <= TXER_IDLE;
                    end if;
                end if;

        end case;
    end process;

    in_o <= accept(config_c, r.state /= ST_SEND_STATS_NO_EOP and 
                             r.state /= ST_SEND_STATS_EOP and 
                             r.state /= ST_REALIGN_BUF and 
                             r.state /= ST_HEADER_STATS and 
                             r.state /= ST_RESET_STATS);

    proc_txer: process(r, in_i)
    begin
        out_o <= transfer_defaults(config_c);
        case r.txer is 
            when TXER_SEND_STATS => 
                out_o <= transfer(config_c,
                                  src => next_beat(stats_buf_config, r.stats_buf, last => false),
                                  force_last => true,
                                  last => is_last(stats_buf_config, r.stats_buf));  
            when others => 
        end case;
    end process;

    assert_proc: process(r,in_i, clock_i)
        variable header_buf, next_header : header_t;
        variable next_header_byte_string,header_byte_sring : byte_string(0 to HEADER_SIZE-1);
    begin 

        header_buf := header_unpack(bytes(header_config_c,r.header_buf), to_integer(r.rx_bytes));

        next_header_byte_string := bytes(header_config_c,shift(header_config_c, r.header_buf, in_i));
        header_byte_sring := bytes(header_config_c,r.header_buf);

        case r.state is

            when ST_HEADER_DEC => 
           

            when ST_HEADER_STATS | ST_REALIGN_BUF =>
                assert to_integer(r.header.pkt_size) <= mtu_c report "ERROR: Size cannot be supp to mtu" severity failure;



            when ST_SEND_STATS_EOP => 
                -- assert r.stats.stats_header_valid and r.stats.stats_payload_valid
                -- report "Error detected"
                -- severity WARNING;

            when others =>

        end case;
    end process;

end architecture;
