  constant SWD_AP_INTERVAL     : std_ulogic_vector(7 downto 0):= "10------";
  constant SWD_AP_ID_HIGH      : std_ulogic_vector(7 downto 0):= "1100----";
  constant SWD_AP_ID_LOW       : std_ulogic_vector(7 downto 0):= "1101----";
  constant SWD_AP_TARGET_ADDR  : std_ulogic_vector(7 downto 0):= "1110----";
  constant SWD_AP_ABORT        : std_ulogic_vector(7 downto 0):= "1111----";
  constant SWD_AP_RW           : std_ulogic_vector(7 downto 0):= "0-------";
  constant SWD_AP_READ         : std_ulogic_vector(7 downto 0):= "00------";
  constant SWD_AP_WRITE        : std_ulogic_vector(7 downto 0):= "01------";
  
