library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library nsl_data, nsl_amba, nsl_math, nsl_logic;
use nsl_data.bytestream.all;
use nsl_amba.axi4_stream.all;
use nsl_data.crc.all;
use nsl_data.prbs.all;
use nsl_amba.random_pkt_checker.all;
use nsl_data.endian.all;

entity random_pkt_generator is
  generic (
    mtu_c: integer := 1500;
    config_c: config_t;
    data_prbs_init_c: prbs_state := x"deadbee"&"111";
    data_prbs_poly_c: prbs_state := prbs31
    );
  port (
    clock_i : in std_ulogic;
    reset_n_i : in std_ulogic;
    --
    in_i : in master_t;
    in_o : out slave_t;
    --
    out_o : out master_t;
    out_i : in slave_t
    );
end entity;

architecture beh of random_pkt_generator is

    constant header_size : integer := 8;
    constant header_config_c : buffer_config_t := buffer_config(config_c, header_size);
    constant cmd_buf_config : buffer_config_t := buffer_config(config_c, cmd_packed_t'length);
    constant mtu_l2 : integer := nsl_math.arith.log2(mtu_c) + 1;
    constant data_width_l2 : integer := nsl_math.arith.log2(config_c.data_width);

    type state_t is (
        ST_RESET,
        ST_CMD_GET,
        ST_CMD_DEC,
        ST_BUILD_HEADER,
        ST_SEND_HEADER,
        ST_SEND_PAYLOAD
        );

    function keep_generator(config_c: config_t; data_remainder : integer; is_last_word : boolean) return std_ulogic_vector is
        variable ret : std_ulogic_vector(0 to config_c.data_width-1) := (others => '1');
    begin 
        if is_last_word then
            if data_remainder /= 0 then
                ret(data_remainder to ret'right) := (others => '0');
            end if;
        end if;
        return ret;
    end function;

    type regs_t is
        record
            state : state_t;
            state_pkt_gen : prbs_state(30 downto 0);
            cmd: cmd_t;
            header : buffer_t;
            cmd_buf : buffer_t;
            data_remainder : integer range 0 to config_c.data_width - 1;
            tx_bytes : unsigned(mtu_l2 - 1 downto 0);
            pkt_has_data : boolean;
        end record;
      
        signal r, rin: regs_t;
begin

    regs: process(reset_n_i, clock_i) is
    begin
      if rising_edge(clock_i) then
        r <= rin;
      end if;
      if reset_n_i = '0' then
        r.state <= ST_RESET;
      end if;
    end process;

    gen_process: process(r, in_i, out_i)
        variable cmd_v : cmd_t;
        variable cmd_byte_v : cmd_packed_t;
    begin

        rin <= r;

        cmd_byte_v := bytes(cmd_buf_config, r.cmd_buf);
        cmd_v := cmd_unpack(cmd_byte_v);

        case r.state is
            when ST_RESET =>
                rin.state <= ST_CMD_GET;
                rin.tx_bytes <= to_unsigned(config_c.data_width, r.tx_bytes'length);
                rin.cmd_buf <= reset(cmd_buf_config);

            when ST_CMD_GET =>
                if is_valid(config_c, in_i) then
                    rin.cmd_buf <= shift(cmd_buf_config, r.cmd_buf, in_i);
                    if is_last(cmd_buf_config, r.cmd_buf) then
                        rin.state <= ST_CMD_DEC;
                    end if;
                end if;

            when ST_CMD_DEC => 
                rin.tx_bytes <= to_unsigned(config_c.data_width, r.tx_bytes'length);
                rin.state_pkt_gen <= prbs_forward(data_prbs_init_c, data_prbs_poly_c,
                                                  std_ulogic_vector(from_le(cmd_byte_v)));
                rin.cmd <= cmd_v;
                rin.data_remainder <= to_integer(cmd_v.pkt_size(data_width_l2 -1 downto 0));
                rin.pkt_has_data <= (cmd_v.pkt_size > header_packed_t'length);
                rin.state <= ST_BUILD_HEADER;

            when ST_BUILD_HEADER => 
                rin.header <= reset(header_config_c, 
                                    header_pack(header_from_cmd(r.cmd)));
                rin.state <= ST_SEND_HEADER;
                                              
            when ST_SEND_HEADER =>   
                if is_ready(config_c, out_i) then
                    rin.tx_bytes <= r.tx_bytes + config_c.data_width;
                    rin.header <= shift(header_config_c, r.header);
                    
                    if is_last(header_config_c, r.header) or r.tx_bytes >= r.cmd.pkt_size then
                        if r.pkt_has_data then 
                            rin.pkt_has_data <= false;
                            rin.state <= ST_SEND_PAYLOAD;
                        else
                            rin.state <= ST_CMD_GET;
                        end if;
                    end if;
                end if;

            when ST_SEND_PAYLOAD => 
                if is_ready(config_c, out_i) then
                    rin.tx_bytes <= r.tx_bytes + config_c.data_width;

                    rin.state_pkt_gen <= prbs_forward(r.state_pkt_gen, 
                                                      data_prbs_poly_c,
                                                      config_c.data_width * 8);
                    if r.tx_bytes >= r.cmd.pkt_size then
                        rin.state <= ST_CMD_GET;
                    end if;
                end if;

            when others => 
                null;
        end case;
    end process;

    proc_txer: process(r)
        variable payload_byte_v : byte_string(0 to config_c.data_width -1);
        variable is_last_word : boolean := false;
    begin

        is_last_word := (is_last(header_config_c, r.header) and
                        r.cmd.pkt_size <= header_packed_t'length) or (r.tx_bytes >= r.cmd.pkt_size);

        out_o <= transfer_defaults(config_c);

        payload_byte_v :=   prbs_byte_string(
                                r.state_pkt_gen, 
                                data_prbs_poly_c, 
                                config_c.data_width);

        case r.state is
            when ST_SEND_HEADER => 
                out_o <=  transfer(config_c,
                                  bytes => r.header.data(0 to config_c.data_width-1),
                                  keep => keep_generator(config_c, r.data_remainder, is_last_word),
                                  valid => true,
                                  last => is_last_word);
                                
            when ST_SEND_PAYLOAD => 
                out_o <= transfer(config_c,
                                  bytes => payload_byte_v,
                                  keep => keep_generator(config_c, r.data_remainder, is_last_word),
                                  last => is_last_word);

            when others =>
        end case;
    end process;
    
    in_o <=  accept(config_c, r.state = ST_CMD_GET);

end architecture;
