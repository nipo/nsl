library ieee;
use ieee.std_logic_1164.all;

entity synth_log is
  generic(
    message_c: string
    );
  port(
    unused_i : in std_ulogic
    );
end entity;

architecture beh of synth_log is

begin

end architecture;
