library ieee;
use ieee.std_logic_1164.all;

entity tb is
end tb;

architecture arch of tb is

  
begin
  
end;
